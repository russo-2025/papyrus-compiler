module main

import time
import os
import pref

import papyrus.ast
import papyrus.parser
import papyrus.checker
import gen.gen_pex
import papyrus.vm
import arrays

const prefs = pref.Preferences {
		paths: []string{}
		mode: .compile
		backend: .pex
		no_cache: true
	}
	
fn vm_run() {
		src_file := 'Scriptname ABCD 
Float Function Sum(int n1, float n2, float n3) global
return (n1 + n2 as int + n3 as int) as float 
EndFunction

Int Function PexInstructionTest(int n1, int n2) global
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0))
	return Sum(11, 12 as Float, Sum(10, 20 as Float, 30.0)) as int
EndFunction'

	mut table := ast.new_table()
	mut global_scope := &ast.Scope{}
	mut ast_file := parser.parse_text("::gen_test.v/src::", src_file, mut table, prefs, mut global_scope)
	mut c := checker.new_checker(table, prefs)
	c.check(mut ast_file)
	assert c.errors.len == 0
	mut pex_file := gen_pex.gen_pex_file(mut ast_file, mut table, prefs)
	
	os.write_file("M:\\_projects_skyrim\\papyrus-compiler\\modules\\tests\\disasm.txt", pex_file.str()) or { panic(err) }

	//func := pex_file.get_function_from_empty_state("ABCD", "PexInstructionTest") or { panic("func not found") }

	mut ctx := vm.create_context()
	ctx.load_pex_file(pex_file)

	mut swa := []f32{}
	mut res := f32(0)
	for _ in 0..135 {
		mut sw := time.new_stopwatch()
		sw.start()
		vres := ctx.call_static("ABCD", "PexInstructionTest", [ vm.create_value_data[i32](22), vm.create_value_data[i32](23)]) or {
			assert false
			panic("err")
		}
		res = vres.get[i32]()
		ms := f32(sw.elapsed().microseconds()) / 1000
		swa << ms
	}

	swa.sort(a < b)
	println(swa)

	swa = swa[3..swa.len-6].clone()
	println(swa)
	ms := arrays.sum(swa) or { f32(-1) } / f32(swa.len)
	assert res == 83

	instr_in_ms := i64(f64(ctx.get_executed_instructions_count())/f64(ms))
	println('end run ${ms} ms; result: ${res}; ${instr_in_ms} instructions/ms')

	//println("res ${res.get[i32]()}")
}

fn main() {
	mut sw := time.new_stopwatch()
	sw.start()

	vm_run()

	ms := f32(sw.elapsed().microseconds()) / 1000
	println('finish $ms ms')
}