module tests
/*
"Scriptname TestSelectiveLoading

Float Function main(Float value, ObjectReference ref)
    ref.GetDisplayName() ; ObjectReference
    ref.GetFormID() ; ObjectReference
    Game.GetPlayer()
  Return value
EndFunction"
*/