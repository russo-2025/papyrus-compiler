module vm